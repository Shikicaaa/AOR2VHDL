library ieee;
	use ieee.std_logic_1164.all;
	use ieee.numeric_std.all;

entity tb is
	generic( n : integer := 4);
end tb;

architecture a_tb of tb is
	signal clk, reset : std_logic;
	signal dout : std_logic_vector(0 to n-1);
begin
	dut: entity work.brojac(a_brojac)
		port map(reset, clk, dout);
	clock: process
	begin
		clk <= '0';
		wait for 50 ns;
		clk <= '1';
		wait for 50 ns;
	end process clock;
	stimulus: process
	begin 
		reset <= '1';
		wait for 350 ns;
		reset <= '0';
		wait for 1 us;
	end process stimulus;
end architecture;